
# 
VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
 TIME NANOSECONDS 1 ;
 CAPACITANCE PICOFARADS 1 ;
 RESISTANCE OHMS 1 ;
 DATABASE MICRONS 1000 ;
END UNITS

MANUFACTURINGGRID 0.005 ;
LAYER GC
 TYPE MASTERSLICE ;
END GC

LAYER M1
 TYPE ROUTING ;
 PITCH 0.56 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.23 ;
 SPACING 0.23 ;
 SPACING 0.23 RANGE 0 9.995 ;
 SPACING 0.6 RANGE 10 100000 ;
 RESISTANCE RPERSQ 0.08 ;
 CAPACITANCE CPERSQDIST 3.51e-05 ;
 AREA 0.202 ;
 MINWIDTH 0.23 ;
 ANTENNASIDEAREARATIO 400 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.203 400 ) ( 0.203001 2281.2 ) ( 1.203 2681.2 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
 THICKNESS 0.54 ;
 HEIGHT 1.05 ;
END M1

LAYER V2
 TYPE CUT ;
 SPACING 0.26 ;
 ANTENNAAREARATIO 20 ;
 ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.203 20 ) ( 0.203001 91.9161 ) ( 1.203 175.246 ) ) ;
 ANTENNAAREAFACTOR 1 ;
END V2

LAYER M2
 TYPE ROUTING ;
 PITCH 0.56 ;
 DIRECTION VERTICAL ;
 WIDTH 0.28 ;
 SPACING 0.28 ;
 SPACING 0.28 RANGE 0 9.995 ;
 SPACING 0.6 RANGE 10 100000 ;
 RESISTANCE RPERSQ 0.08 ;
 CAPACITANCE CPERSQDIST 1.46e-05 ;
 AREA 0.202 ;
 MINWIDTH 0.28 ;
 ANTENNASIDEAREARATIO 400 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.203 400 ) ( 0.203001 2281.2 ) ( 1.203 2681.2 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
 THICKNESS 0.54 ;
 HEIGHT 2.41 ;
END M2

LAYER V3
 TYPE CUT ;
 SPACING 0.26 ;
 ANTENNAAREARATIO 20 ;
 ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.203 20 ) ( 0.203001 91.9161 ) ( 1.203 175.246 ) ) ;
 ANTENNAAREAFACTOR 1 ;
END V3

LAYER M3
 TYPE ROUTING ;
 PITCH 0.84 ;
 DIRECTION HORIZONTAL ;
 WIDTH 0.28 ;
 SPACING 0.28 ;
 SPACING 0.28 RANGE 0 9.995 ;
 SPACING 0.6 RANGE 10 100000 ;
 RESISTANCE RPERSQ 0.08 ;
 CAPACITANCE CPERSQDIST 9.24e-06 ;
 AREA 0.202 ;
 MINWIDTH 0.28 ;
 ANTENNASIDEAREARATIO 400 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.203 400 ) ( 0.203001 2281.2 ) ( 1.203 2681.2 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
 THICKNESS 0.54 ;
 HEIGHT 3.77 ;
END M3

LAYER TOP_V
 TYPE CUT ;
 SPACING 0.35 ;
 ANTENNAAREARATIO 20 ;
 ANTENNADIFFAREARATIO PWL ( ( 0 20 ) ( 0.203 20 ) ( 0.203001 91.9161 ) ( 1.203 175.246 ) ) ;
 ANTENNAAREAFACTOR 1 ;
END TOP_V

LAYER TOP_M
 TYPE ROUTING ;
 PITCH 1.12 ;
 DIRECTION VERTICAL ;
 WIDTH 0.44 ;
 SPACING 0.46 ;
 SPACING 0.46 RANGE 0 9.995 ;
 SPACING 0.6 RANGE 10 100000 ;
 RESISTANCE RPERSQ 0.04 ;
 CAPACITANCE CPERSQDIST 4.389e-06 ;
 AREA 0.562 ;
 MINWIDTH 0.44 ;
 ANTENNASIDEAREARATIO 400 ;
 ANTENNADIFFSIDEAREARATIO PWL ( ( 0 400 ) ( 0.203 400 ) ( 0.203001 31624 ) ( 1.203 39624 ) ) ;
 ANTENNASIDEAREAFACTOR 1 ;
 THICKNESS 0.84 ;
 HEIGHT 5.11 ;
END TOP_M

LAYER OverlapCheck
 TYPE OVERLAP ;
END OverlapCheck


VIA V2 DEFAULT
LAYER M1 ;
 RECT -0.14 -0.19 0.14 0.19 ;
LAYER V2 ;
 RECT -0.13 -0.13 0.13 0.13 ;
LAYER M2 ;
 RECT -0.14 -0.19 0.14 0.19 ;
 RESISTANCE 6 ;
END V2

VIA V3 DEFAULT
LAYER M2 ;
 RECT -0.19 -0.14 0.19 0.14 ;
LAYER V3 ;
 RECT -0.13 -0.13 0.13 0.13 ;
LAYER M3 ;
 RECT -0.19 -0.14 0.19 0.14 ;

 RESISTANCE 6 ;
END V3

VIA VL DEFAULT
LAYER M3 ;
 RECT -0.19 -0.24 0.19 0.24 ;
LAYER TOP_V ;
 RECT -0.18 -0.18 0.18 0.18 ;
LAYER TOP_M ;
 RECT -0.27 -0.27 0.27 0.27 ;

 RESISTANCE 2.5 ;
END VL

VIA V2_cross DEFAULT
LAYER M1 ;
 RECT -0.19 -0.14 0.19 0.14 ;
LAYER V2 ;
 RECT -0.13 -0.13 0.13 0.13 ;
LAYER M2 ;
 RECT -0.14 -0.19 0.14 0.19 ;

 RESISTANCE 6 ;
END V2_cross

VIA V3_cross DEFAULT
LAYER M2 ;
 RECT -0.14 -0.19 0.14 0.19 ;
LAYER V3 ;
 RECT -0.13 -0.13 0.13 0.13 ;
LAYER M3 ;
 RECT -0.19 -0.14 0.19 0.14 ;

 RESISTANCE 6 ;
END V3_cross


VIA V3_TOS_N DEFAULT TOPOFSTACKONLY
RESISTANCE 6.00 ;
LAYER M2 ;
    RECT -0.14 -0.19 0.14 0.535 ;
LAYER V3 ;
    RECT -0.13 -0.13 0.13 0.13 ;
LAYER M3 ;
    RECT -0.19 -0.14 0.19 0.14 ;
END V3_TOS_N

VIA V3_TOS_S DEFAULT TOPOFSTACKONLY
RESISTANCE 6.00 ;
LAYER M2 ;
    RECT -0.14 -0.535 0.14 0.19 ;
LAYER V3 ;
    RECT -0.13 -0.13 0.13 0.13 ;
LAYER M3 ;
    RECT -0.19 -0.14 0.19 0.14 ;
END V3_TOS_S

VIA VL_TOS_E DEFAULT TOPOFSTACKONLY
RESISTANCE 2.5 ;
LAYER M3 ;
    RECT -0.24 -0.19 0.485 0.19 ;
LAYER TOP_V ;
    RECT -0.18 -0.18 0.18 0.18 ;
LAYER TOP_M ;
    RECT -0.27 -0.27 0.27 0.27 ;
END VL_TOS_E

VIA VL_TOS_W DEFAULT TOPOFSTACKONLY
RESISTANCE 2.5 ;
LAYER M3 ;
    RECT -0.485 -0.19 0.24 0.19 ;
LAYER TOP_V ;
    RECT -0.18 -0.18 0.18 0.18 ;
LAYER TOP_M ;
    RECT -0.27 -0.27 0.27 0.27 ;
END VL_TOS_W


VIARULE V2 GENERATE
    LAYER M1 ;
 	ENCLOSURE 0.06 0.01 ;
    LAYER M2 ;
 	ENCLOSURE 0.06 0.01 ;
    LAYER V2 ;
        RECT -0.13 -0.13 0.13 0.13 ;
        SPACING 0.52 BY 0.52 ;
END V2

VIARULE V3 GENERATE
    LAYER M2 ;
 	ENCLOSURE 0.06 0.01 ;
    LAYER M3 ;
 	ENCLOSURE 0.06 0.01 ;
    LAYER V3 ;
        RECT -0.13 -0.13 0.13 0.13 ;
        SPACING 0.52 BY 0.52 ;
END V3

VIARULE VL GENERATE
    LAYER M3 ;
 	ENCLOSURE 0.06 0.01 ;
    LAYER TOP_M ;
 	ENCLOSURE 0.09 0.09 ;
    LAYER TOP_V ;
        RECT -0.18 -0.18 0.18 0.18 ;
        SPACING 0.71 BY 0.71 ;
END VL

END LIBRARY
